module pattern_table(addr, data, out, mode);
	input wire[10:0] addr;
	input wire[1:0] data;
	input wire mode;
	output reg[1:0] out;
	
endmodule
module ricardo (a,b);

input a;
output reg b;

endmodule 